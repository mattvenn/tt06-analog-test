magic
tech sky130A
magscale 1 2
timestamp 1707993328
<< pwell >>
rect -201 -7534 201 7534
<< psubdiff >>
rect -165 7464 -69 7498
rect 69 7464 165 7498
rect -165 7402 -131 7464
rect 131 7402 165 7464
rect -165 -7464 -131 -7402
rect 131 -7464 165 -7402
rect -165 -7498 -69 -7464
rect 69 -7498 165 -7464
<< psubdiffcont >>
rect -69 7464 69 7498
rect -165 -7402 -131 7402
rect 131 -7402 165 7402
rect -69 -7498 69 -7464
<< xpolycontact >>
rect -35 6936 35 7368
rect -35 4504 35 4936
rect -35 3968 35 4400
rect -35 1536 35 1968
rect -35 1000 35 1432
rect -35 -1432 35 -1000
rect -35 -1968 35 -1536
rect -35 -4400 35 -3968
rect -35 -4936 35 -4504
rect -35 -7368 35 -6936
<< ppolyres >>
rect -35 4936 35 6936
rect -35 1968 35 3968
rect -35 -1000 35 1000
rect -35 -3968 35 -1968
rect -35 -6936 35 -4936
<< locali >>
rect -165 7464 -69 7498
rect 69 7464 165 7498
rect -165 7402 -131 7464
rect 131 7402 165 7464
rect -165 -7464 -131 -7402
rect 131 -7464 165 -7402
rect -165 -7498 -69 -7464
rect 69 -7498 165 -7464
<< viali >>
rect -19 6953 19 7350
rect -19 4522 19 4919
rect -19 3985 19 4382
rect -19 1554 19 1951
rect -19 1017 19 1414
rect -19 -1414 19 -1017
rect -19 -1951 19 -1554
rect -19 -4382 19 -3985
rect -19 -4919 19 -4522
rect -19 -7350 19 -6953
<< metal1 >>
rect -25 7350 25 7362
rect -25 6953 -19 7350
rect 19 6953 25 7350
rect -25 6941 25 6953
rect -25 4919 25 4931
rect -25 4522 -19 4919
rect 19 4522 25 4919
rect -25 4510 25 4522
rect -25 4382 25 4394
rect -25 3985 -19 4382
rect 19 3985 25 4382
rect -25 3973 25 3985
rect -25 1951 25 1963
rect -25 1554 -19 1951
rect 19 1554 25 1951
rect -25 1542 25 1554
rect -25 1414 25 1426
rect -25 1017 -19 1414
rect 19 1017 25 1414
rect -25 1005 25 1017
rect -25 -1017 25 -1005
rect -25 -1414 -19 -1017
rect 19 -1414 25 -1017
rect -25 -1426 25 -1414
rect -25 -1554 25 -1542
rect -25 -1951 -19 -1554
rect 19 -1951 25 -1554
rect -25 -1963 25 -1951
rect -25 -3985 25 -3973
rect -25 -4382 -19 -3985
rect 19 -4382 25 -3985
rect -25 -4394 25 -4382
rect -25 -4522 25 -4510
rect -25 -4919 -19 -4522
rect 19 -4919 25 -4522
rect -25 -4931 25 -4919
rect -25 -6953 25 -6941
rect -25 -7350 -19 -6953
rect 19 -7350 25 -6953
rect -25 -7362 25 -7350
<< properties >>
string FIXED_BBOX -148 -7481 148 7481
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.35 l 10.0 m 5 nx 1 wmin 0.350 lmin 0.50 rho 319.8 val 10.25k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
