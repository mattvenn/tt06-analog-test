magic
tech sky130A
magscale 1 2
timestamp 1707991876
<< metal1 >>
rect 18398 42349 23025 42882
rect 18398 41873 18931 42349
rect 18398 41656 20410 41873
rect 18398 41340 20440 41656
rect 20060 41136 20440 41340
rect 20494 41606 20998 41658
rect 20494 41554 21472 41606
rect 20494 41378 21654 41554
rect 20494 41100 21472 41378
rect 9692 40716 9702 40748
rect 9518 40364 9702 40716
rect 9692 40132 9702 40364
rect 10302 40716 10312 40748
rect 10302 40686 20032 40716
rect 20950 40686 21472 41100
rect 10302 40460 21472 40686
rect 10302 40364 20032 40460
rect 10302 40132 10312 40364
rect 20950 3202 21472 40460
rect 22492 4855 23025 42349
rect 31066 4855 31602 4856
rect 22492 4322 31602 4855
rect 20950 2680 27071 3202
rect 26549 1964 27071 2680
rect 31066 2000 31602 4322
rect 26512 1216 26522 1964
rect 27362 1216 27372 1964
rect 31006 1400 31016 2000
rect 31642 1400 31652 2000
<< via1 >>
rect 9702 40132 10302 40748
rect 26522 1216 27362 1964
rect 31016 1400 31642 2000
<< metal2 >>
rect 9702 40748 10302 40758
rect 9702 40122 10302 40132
rect 31016 2000 31642 2010
rect 26522 1964 27362 1974
rect 31016 1390 31642 1400
rect 26522 1206 27362 1216
<< via2 >>
rect 9702 40132 10302 40748
rect 26522 1216 27362 1964
rect 31016 1400 31642 2000
<< metal3 >>
rect 9692 40748 10312 40753
rect 9692 40132 9702 40748
rect 10302 40132 10312 40748
rect 9692 40127 10312 40132
rect 31006 2000 31652 2005
rect 26512 1964 27372 1969
rect 26512 1216 26522 1964
rect 27362 1216 27372 1964
rect 31006 1400 31016 2000
rect 31642 1400 31652 2000
rect 31006 1395 31652 1400
rect 26512 1211 27372 1216
<< via3 >>
rect 9702 40132 10302 40748
rect 26522 1216 27362 1964
rect 31016 1400 31642 2000
<< metal4 >>
rect 200 200 500 45152
rect 798 44952 858 45152
rect 1534 44952 1594 45152
rect 2270 44952 2330 45152
rect 3006 44952 3066 45152
rect 3742 44952 3802 45152
rect 4478 44952 4538 45152
rect 5214 44952 5274 45152
rect 5950 44952 6010 45152
rect 6686 44952 6746 45152
rect 7422 44952 7482 45152
rect 8158 44952 8218 45152
rect 8894 44952 8954 45152
rect 9630 44952 9690 45152
rect 9800 40749 10100 45152
rect 10366 44952 10426 45152
rect 11102 44952 11162 45152
rect 11838 44952 11898 45152
rect 12574 44952 12634 45152
rect 13310 44952 13370 45152
rect 14046 44952 14106 45152
rect 14782 44952 14842 45152
rect 15518 44952 15578 45152
rect 16254 44952 16314 45152
rect 16990 44952 17050 45152
rect 17726 44952 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44952 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 9701 40748 10303 40749
rect 9701 40132 9702 40748
rect 10302 40132 10303 40748
rect 9701 40131 10303 40132
rect 200 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 200
rect 9800 0 10100 40131
rect 31015 2000 31643 2001
rect 26521 1964 27363 1965
rect 26521 1216 26522 1964
rect 27362 1216 27363 1964
rect 31015 1400 31016 2000
rect 31642 1400 31643 2000
rect 31015 1399 31643 1400
rect 26521 1215 27363 1216
rect 26836 200 27014 1215
rect 13648 0 13768 200
rect 18064 0 18184 200
rect 22480 0 22600 200
rect 26836 0 27016 200
rect 26836 -8 27014 0
rect 31296 -34 31474 1399
<< via4 >>
rect 9702 40132 10302 40748
rect 26522 1216 27362 1964
rect 31016 1400 31642 2000
<< metal5 >>
rect 9678 40748 10326 40772
rect 9678 40132 9702 40748
rect 10302 40132 10326 40748
rect 9678 40108 10326 40132
rect 30992 2000 31666 2024
rect 26498 1964 27386 1988
rect 26498 1216 26522 1964
rect 27362 1216 27386 1964
rect 30992 1400 31016 2000
rect 31642 1400 31666 2000
rect 30992 1376 31666 1400
rect 26498 1192 27386 1216
use sky130_fd_pr__res_high_po_0p35_EB2D9Q  sky130_fd_pr__res_high_po_0p35_EB2D9Q_0
timestamp 1707991876
transform 1 0 20533 0 1 40898
box -367 -482 367 482
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal tristate
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal tristate
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal tristate
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal tristate
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal tristate
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal tristate
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal tristate
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal tristate
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal tristate
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal tristate
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal tristate
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal tristate
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal tristate
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal tristate
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal tristate
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal tristate
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal tristate
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal tristate
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal tristate
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal tristate
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal tristate
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal tristate
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal tristate
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal tristate
flabel metal4 200 0 500 45152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel space 9800 0 10100 45152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
