magic
tech sky130A
magscale 1 2
timestamp 1707993328
<< poly >>
rect -249 579 -183 595
rect -249 545 -233 579
rect -199 545 -183 579
rect -249 165 -183 545
rect -249 -545 -183 -165
rect -249 -579 -233 -545
rect -199 -579 -183 -545
rect -249 -595 -183 -579
rect -141 579 -75 595
rect -141 545 -125 579
rect -91 545 -75 579
rect -141 165 -75 545
rect -141 -545 -75 -165
rect -141 -579 -125 -545
rect -91 -579 -75 -545
rect -141 -595 -75 -579
rect -33 579 33 595
rect -33 545 -17 579
rect 17 545 33 579
rect -33 165 33 545
rect -33 -545 33 -165
rect -33 -579 -17 -545
rect 17 -579 33 -545
rect -33 -595 33 -579
rect 75 579 141 595
rect 75 545 91 579
rect 125 545 141 579
rect 75 165 141 545
rect 75 -545 141 -165
rect 75 -579 91 -545
rect 125 -579 141 -545
rect 75 -595 141 -579
rect 183 579 249 595
rect 183 545 199 579
rect 233 545 249 579
rect 183 165 249 545
rect 183 -545 249 -165
rect 183 -579 199 -545
rect 233 -579 249 -545
rect 183 -595 249 -579
<< polycont >>
rect -233 545 -199 579
rect -233 -579 -199 -545
rect -125 545 -91 579
rect -125 -579 -91 -545
rect -17 545 17 579
rect -17 -579 17 -545
rect 91 545 125 579
rect 91 -579 125 -545
rect 199 545 233 579
rect 199 -579 233 -545
<< npolyres >>
rect -249 -165 -183 165
rect -141 -165 -75 165
rect -33 -165 33 165
rect 75 -165 141 165
rect 183 -165 249 165
<< locali >>
rect -249 545 -233 579
rect -199 545 -183 579
rect -141 545 -125 579
rect -91 545 -75 579
rect -33 545 -17 579
rect 17 545 33 579
rect 75 545 91 579
rect 125 545 141 579
rect 183 545 199 579
rect 233 545 249 579
rect -249 -579 -233 -545
rect -199 -579 -183 -545
rect -141 -579 -125 -545
rect -91 -579 -75 -545
rect -33 -579 -17 -545
rect 17 -579 33 -545
rect 75 -579 91 -545
rect 125 -579 141 -545
rect 183 -579 199 -545
rect 233 -579 249 -545
<< viali >>
rect -233 545 -199 579
rect -125 545 -91 579
rect -17 545 17 579
rect 91 545 125 579
rect 199 545 233 579
rect -233 182 -199 545
rect -125 182 -91 545
rect -17 182 17 545
rect 91 182 125 545
rect 199 182 233 545
rect -233 -545 -199 -182
rect -125 -545 -91 -182
rect -17 -545 17 -182
rect 91 -545 125 -182
rect 199 -545 233 -182
rect -233 -579 -199 -545
rect -125 -579 -91 -545
rect -17 -579 17 -545
rect 91 -579 125 -545
rect 199 -579 233 -545
<< metal1 >>
rect -239 579 -193 591
rect -239 182 -233 579
rect -199 182 -193 579
rect -239 170 -193 182
rect -131 579 -85 591
rect -131 182 -125 579
rect -91 182 -85 579
rect -131 170 -85 182
rect -23 579 23 591
rect -23 182 -17 579
rect 17 182 23 579
rect -23 170 23 182
rect 85 579 131 591
rect 85 182 91 579
rect 125 182 131 579
rect 85 170 131 182
rect 193 579 239 591
rect 193 182 199 579
rect 233 182 239 579
rect 193 170 239 182
rect -239 -182 -193 -170
rect -239 -579 -233 -182
rect -199 -579 -193 -182
rect -239 -591 -193 -579
rect -131 -182 -85 -170
rect -131 -579 -125 -182
rect -91 -579 -85 -182
rect -131 -591 -85 -579
rect -23 -182 23 -170
rect -23 -579 -17 -182
rect 17 -579 23 -182
rect -23 -591 23 -579
rect 85 -182 131 -170
rect 85 -579 91 -182
rect 125 -579 131 -182
rect 85 -591 131 -579
rect 193 -182 239 -170
rect 193 -579 199 -182
rect 233 -579 239 -182
rect 193 -591 239 -579
<< properties >>
string gencell sky130_fd_pr__res_generic_po
string library sky130
string parameters w 0.33 l 1.65 m 1 nx 5 wmin 0.330 lmin 1.650 rho 48.2 val 241.0 dummy 0 dw 0.0 term 0.0 sterm 0.0 caplen 0.4 snake 0 guard 0 glc 1 grc 1 gtc 1 gbc 1 roverlap 0 endcov 100 full_metal 1 hv_guard 0 n_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
